
`ifndef RKV_I2C_USER_ELEMENT_SEQUENCES_SVH
`define RKV_I2C_USER_ELEMENT_SEQUENCES_SVH

`include "rkv_apb_user_config_seq.sv"
`include "rkv_user_wait_detect_abort_source_seq.sv"
`include "rkv_i2c_master_abrt_sbyte_norstrt_virt_seq.sv"
`include "rkv_apb_noread_packet_seq.sv"
`include "rkv_apb_write_nocheck_packet_seq.sv"
`endif // RKV_I2C_USER_ELEMENT_SEQUENCES_SVH

 